interface intf;
  logic x;
  logic y;
  logic z;
  logic borrow;
  logic diff;
endinterface
